work.fulladder(main) rtlc_no_parameters
